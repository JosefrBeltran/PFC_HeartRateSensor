** Profile: "SCHEMATIC1-Herat_Rate_Amplifier"  [ C:\Users\josefr\Dropbox\Upct\Proyecto\Design\heart_rate_amplifier-SCHEMATIC1-Herat_Rate_Amplifier.sim ] 

** Creating circuit file "heart_rate_amplifier-SCHEMATIC1-Herat_Rate_Amplifier.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of c:\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 2s 3 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\heart_rate_amplifier-SCHEMATIC1.net" 


.END
